// These pins should all exist in ice40.pcf
input clk_100p0,
// RGB LED
inout ICE_39,
inout ICE_40,
inout ICE_41,
// UART
inout ICE_25,
inout ICE_27,
// PMODs for VGA demo
// PMOD0A
inout ICE_45,
inout ICE_47,
inout ICE_2,
inout ICE_4,
// PMOD0B
inout ICE_44,
inout ICE_46,
inout ICE_48,
inout ICE_3,
// PMOD1A
inout ICE_31,
inout ICE_34,
inout ICE_38,
inout ICE_43,
// PMOD1B
inout ICE_28,
inout ICE_32,
inout ICE_36,
inout ICE_42
